module test (
    reset,
    clk,
    data_i,
    data_o
    );

    input               reset;
    input               clk;
    input [8:0]         data_i;
    output [8:0]        data_o;

endmodule

